module RAM16x59S (WCLK,addr,I,O);
  input WCLK;
  input [3:0] addr;
  input [58:0] I;
  output [58:0] O;
    
  wire WCLK;
  wire [3:0] addr;
  wire [58:0] I;
  wire [58:0] O;

  RAM16X1S #(.INIT(16'h0000)) RAM_0 (.O(O[0]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[0]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_1 (.O(O[1]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[1]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_2 (.O(O[2]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[2]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_3 (.O(O[3]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[3]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_4 (.O(O[4]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[4]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_5 (.O(O[5]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[5]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_6 (.O(O[6]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[6]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_7 (.O(O[7]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[7]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_8 (.O(O[8]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[8]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_9 (.O(O[9]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[9]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_10 (.O(O[10]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[10]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_11 (.O(O[11]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[11]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_12 (.O(O[12]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[12]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_13 (.O(O[13]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[13]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_14 (.O(O[14]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[14]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_15 (.O(O[15]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[15]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_16 (.O(O[16]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[16]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_17 (.O(O[17]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[17]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_18 (.O(O[18]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[18]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_19 (.O(O[19]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[19]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_20 (.O(O[20]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[20]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_21 (.O(O[21]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[21]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_22 (.O(O[22]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[22]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_23 (.O(O[23]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[23]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_24 (.O(O[24]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[24]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_25 (.O(O[25]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[25]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_26 (.O(O[26]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[26]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_27 (.O(O[27]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[27]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_28 (.O(O[28]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[28]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_29 (.O(O[29]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[29]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_30 (.O(O[30]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[30]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_31 (.O(O[31]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[31]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_32 (.O(O[32]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[32]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_33 (.O(O[33]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[33]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_34 (.O(O[34]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[34]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_35 (.O(O[35]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[35]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_36 (.O(O[36]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[36]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_37 (.O(O[37]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[37]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_38 (.O(O[38]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[38]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_39 (.O(O[39]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[39]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_40 (.O(O[40]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[40]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_41 (.O(O[41]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[41]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_42 (.O(O[42]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[42]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_43 (.O(O[43]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[43]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_44 (.O(O[44]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[44]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_45 (.O(O[45]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[45]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_46 (.O(O[46]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[46]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_47 (.O(O[47]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[47]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_48 (.O(O[48]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[48]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_49 (.O(O[49]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[49]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_50 (.O(O[50]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[50]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_51 (.O(O[51]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[51]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_52 (.O(O[52]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[52]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_53 (.O(O[53]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[53]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_54 (.O(O[54]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[54]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_55 (.O(O[55]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[55]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_56 (.O(O[56]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[56]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_57 (.O(O[57]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[57]),.WCLK(WCLK),.WE(1'b1));
  RAM16X1S #(.INIT(16'h0000)) RAM_58 (.O(O[58]),.A0(addr[0]),.A1(addr[1]),.A2(addr[2]),.A3(addr[3]),.D(I[58]),.WCLK(WCLK),.WE(1'b1));
endmodule

