// THIS FILE HAS BEEN MODIFIED BY fixpsmV (Scott Gravenhorst)
// Comments delimited by /* and */ have been removed.

`timescale 1 ps / 1ps
module midictrl (address, instruction, proc_reset, clk);
input  [9:0]  address;
input   clk ;
output  [17:0]  instruction ;
output   proc_reset ;
wire  [10:0] jaddr ;
wire  [0:0] jparity ;
wire   [7:0] jdata ;
wire   [7:0] doa ;
wire   [0:0] dopa ;
wire   tdo1 ;
wire   tdo2 ;
wire   update ;
wire   shift  ;
wire   reset  ;
wire   tdi  ;
wire   sel1 ;
wire   drck1  ;
wire   drck1_buf ;
wire   sel2 ;
wire   drck2  ;
wire   capture ;
wire   tap5 ;
wire   tap11  ;
wire   tap17  ;
RAMB16_S9_S18 ram_1024_x_18(
 .DIB  (16'h0000),
 .DIPB  (2'b00),
 .ENB (1'b1),
 .WEB (1'b0),
 .SSRB (1'b0),
 .CLKB (clk),
 .ADDRB (address),
 .DOB (instruction[15:0]),
 .DOPB (instruction[17:16]),
 .DIA  (jdata),
 .DIPA  (jparity),
 .ENA (sel1),
 .WEA (1'b1),
 .SSRA (1'b0),
 .CLKA (update),
 .ADDRA (jaddr),
 .DOA (doa[7:0]),
 .DOPA (dopa))
;
defparam ram_1024_x_18.INIT_00  = 256'hCFF6CFF2CFF9CFF80F000B000800070006000500040001000A000000C2FF00E9;
defparam ram_1024_x_18.INIT_01  = 256'h603E4021AAFD603F50162A02541F2A0154802A04C001EF000FFFCFF10F40EF3D;
defparam ram_1024_x_18.INIT_02  = 256'h4B0550454B0450404B03503B4B0250364B01504F4B0054672080501640FEAAFE;
defparam ram_1024_x_18.INIT_03  = 256'h40160B7F501640000B0340160B7F5016407F0B02401650164B7F504C4B065049;
defparam ram_1024_x_18.INIT_04  = 256'hC4014016D0E00B7F40161E000B064016CEE01E000B0540160B7F501640000B04;
defparam ram_1024_x_18.INIT_05  = 256'h50612F800F005C5E9FE00E0A0E064E071F604016505742805057429016005063;
defparam ram_1024_x_18.INIT_06  = 256'h0B00547140F7547542F0A30FA2F01300120040161450CA041700401616F00F7F;
defparam ram_1024_x_18.INIT_07  = 256'h401615400401407E0402507D42D0507D42C019000B0040160B01541640F04016;
defparam ram_1024_x_18.INIT_08  = 256'h42B050DC42A05098429050A94280A2F01210119054165DF04D02AF0F1F90AAFB;
defparam ram_1024_x_18.INIT_09  = 256'h880150A0483CF680C614C7F950A94700401650D942E050D742D050DC42C050C3;
defparam ram_1024_x_18.INIT_0A  = 256'h7FE00E0050C0C80150C04800C6144016CFF80F01CFF80F0050164700CDFA1D60;
defparam ram_1024_x_18.INIT_0B  = 256'h40A188017D80C80140AF8E0140B38D01FFD07FE08E0150BC5D801DE054BA5F60;
defparam ram_1024_x_18.INIT_0C  = 256'h46114016C7F454CF46104016C7F754CB46404016C7F354C746014016CFF80F00;
defparam ram_1024_x_18.INIT_0D  = 256'h58E2CF0C0E0040164016C6F2C7F14016C7F040C008005416467B4016C7F554D3;
defparam ram_1024_x_18.INIT_0E  = 256'h015C0561015C0557012905100146A000DFE00E060E060E060E068F0C40DE8E01;
defparam ram_1024_x_18.INIT_0F  = 256'h015C0520015C0565015C0564015C0569015C0575015C0547015C0565015C0576;
defparam ram_1024_x_18.INIT_10  = 256'h015C052E015C055301290520015C0568015C0574015C056E015C0579015C0553;
defparam ram_1024_x_18.INIT_11  = 256'h015C0568015C056E015C0565015C0576015C0561015C0572015C0547015C0520;
defparam ram_1024_x_18.INIT_12  = 256'hA50FA0000133C580A50F512F2510A000015C0574015C0573015C0572015C056F;
defparam ram_1024_x_18.INIT_13  = 256'h04F0017701420406040604060407145001730142C408A4F01450A0000133C5C0;
defparam ram_1024_x_18.INIT_14  = 256'h0142042001770142017C01420181014204300181A000016DC490A4F8A000C490;
defparam ram_1024_x_18.INIT_15  = 256'hC490C40CA4F01450A000017C017C013305010133050C01330506013305280177;
defparam ram_1024_x_18.INIT_16  = 256'h0173C490E401A000C49004F00177016DC490040604060407040714500173016D;
defparam ram_1024_x_18.INIT_17  = 256'h557DC20101770219A0005578C10101730128A0005574C001000BA000C490E401;
defparam ram_1024_x_18.INIT_18  = 256'h51932A40DAC0ACC04C00A0005587C40101810432A0005582C301017C0314A000;
defparam ram_1024_x_18.INIT_19  = 256'h0000000000000000000000008001AA3FCA02EC3F4C0851982A80CA01EC3E4C01;
defparam ram_1024_x_18.INIT_1A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_20  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_21  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_22  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_23  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_24  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_25  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_26  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_27  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_28  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_29  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_30  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_31  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_32  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_33  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_34  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_35  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_36  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_37  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_38  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_39  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3F  = 256'h418B000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_00 = 256'hC337433737403030D3683DD378C38334CD334F777777777430DDDE22AA00000B;
defparam ram_1024_x_18.INITP_01 = 256'hCCCCCCCCCCCE2A9DD3EBB37B7B7B7B78D1DD874D0DD788D8766DF77777740D00;
defparam ram_1024_x_18.INITP_02 = 256'hDCB72D28E28FAA8F80BF3333CFFF3B8A3EA8F02C2C36CCCCCCCCCCCCCCCCCCCC;
defparam ram_1024_x_18.INITP_03 = 256'h000000000000000000000000000000000000000000000000000C2348D02DCB72;
defparam ram_1024_x_18.INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_07 = 256'hC000000000000000000000000000000000000000000000000000000000000000;
  BSCAN_SPARTAN3 v2_bscan(   
       .TDO1(tdo1),
       .TDO2(tdo2),
            .UPDATE(update),
             .SHIFT(shift),
             .RESET(reset),
               .TDI(tdi),
              .SEL1(sel1),
             .DRCK1(drck1),
              .SEL2(sel2),
             .DRCK2(drck2),
    .CAPTURE(capture));
    
  //buffer signal used as a clock
  BUFG upload_clock(
          .I(drck1),
          .O(drck1_buf));
  // Assign the reset to be active whenever the uploading subsystem is active
  assign proc_reset = sel1;
  defparam srlC1.INIT = 16'h0000;
  SRLC16E srlC1 (   
              .D(tdi),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[10]),
            .Q15(jaddr[8]));
            
  FD flop1(
             .D(jaddr[10]),
             .Q(jaddr[9]),
             .C(drck1_buf));
  defparam srlC2.INIT = 16'h0000;
  SRLC16E srlC2 (   
              .D(jaddr[8]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[7]),
            .Q15(tap5));
            
  FD flop2 ( 
             .D(jaddr[7]),
             .Q(jaddr[6]),
             .C(drck1_buf));
  defparam srlC3.INIT = 16'h0000;
  SRLC16E srlC3(   
              .D(tap5),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[5]),
            .Q15(jaddr[3]));
  
  FD flop3 ( 
             .D(jaddr[5]),
             .Q(jaddr[4]),
             .C(drck1_buf));
  defparam srlC4.INIT = 16'h0000;
  SRLC16E srlC4 (   
              .D(jaddr[3]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[2]),
            .Q15(tap11));
  
  FD flop4 ( 
             .D(jaddr[2]),
             .Q(jaddr[1]),
             .C(drck1_buf));
  defparam srlC5.INIT = 16'h0000;
  SRLC16E srlC5 (   
              .D(tap11),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[0]),
            .Q15(jdata[7]));
            
  FD flop5 ( 
             .D(jaddr[0]),
             .Q(jparity[0]),
             .C(drck1_buf));
  defparam srlC6.INIT = 16'h0000;
    SRLC16E srlC6(   
             .D(jdata[7]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[6]),
            .Q15(tap17));
  
  FD flop6 ( 
             .D(jdata[6]),
             .Q(jdata[5]),
             .C(drck1_buf));
  defparam srlC7.INIT = 16'h0000;
  SRLC16E srlC7 (   
              .D(tap17),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[4]),
            .Q15(jdata[2]));
  
  FD flop7 ( 
             .D(jdata[4]),
             .Q(jdata[3]),
             .C(drck1_buf));
  defparam srlC8.INIT = 16'h0000;
  SRLC16E srlC8 (   
             .D(jdata[2]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[1]),
            .Q15(tdo1));
  FD flop8 ( 
             .D(jdata[1]),
             .Q(jdata[0]),
             .C(drck1_buf));
endmodule
