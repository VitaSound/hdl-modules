// THIS FILE HAS BEEN MODIFIED BY fixpsmV (Scott Gravenhorst)
// Comments delimited by /* and */ have been removed.

`timescale 1 ps / 1ps
module midictrl (address, instruction, proc_reset, clk);
input  [9:0]  address;
input   clk ;
output  [17:0]  instruction ;
output   proc_reset ;
wire  [10:0] jaddr ;
wire  [0:0] jparity ;
wire   [7:0] jdata ;
wire   [7:0] doa ;
wire   [0:0] dopa ;
wire   tdo1 ;
wire   tdo2 ;
wire   update ;
wire   shift  ;
wire   reset  ;
wire   tdi  ;
wire   sel1 ;
wire   drck1  ;
wire   drck1_buf ;
wire   sel2 ;
wire   drck2  ;
wire   capture ;
wire   tap5 ;
wire   tap11  ;
wire   tap17  ;
RAMB16_S9_S18 ram_1024_x_18(
 .DIB  (16'h0000),
 .DIPB  (2'b00),
 .ENB (1'b1),
 .WEB (1'b0),
 .SSRB (1'b0),
 .CLKB (clk),
 .ADDRB (address),
 .DOB (instruction[15:0]),
 .DOPB (instruction[17:16]),
 .DIA  (jdata),
 .DIPA  (jparity),
 .ENA (sel1),
 .WEA (1'b1),
 .SSRA (1'b0),
 .CLKA (update),
 .ADDRA (jaddr),
 .DOA (doa[7:0]),
 .DOPA (dopa))
;
defparam ram_1024_x_18.INIT_00  = 256'hCFF6CFF2CFF9CFF80F000B000800070006000500040001000A000000C2FF0111;
defparam ram_1024_x_18.INIT_01  = 256'h603E4021AAFD603F50162A02541F2A0154802A04C001EF000FFFCFF10F40EF3D;
defparam ram_1024_x_18.INIT_02  = 256'h4B0550454B0450404B03503B4B0250364B01504F4B0054672080501640FEAAFE;
defparam ram_1024_x_18.INIT_03  = 256'h40160B7F501640000B0340160B7F5016407F0B02401650164B7F504C4B065049;
defparam ram_1024_x_18.INIT_04  = 256'hC4014016D0E00B7F40161E000B064016CEE01E000B0540160B7F501640000B04;
defparam ram_1024_x_18.INIT_05  = 256'h50612F800F005C5E9FE00E0A0E064E071F604016505742805057429016005063;
defparam ram_1024_x_18.INIT_06  = 256'h0B00547140F7547542F0A30FA2F01300120040161450CA041700401616F00F7F;
defparam ram_1024_x_18.INIT_07  = 256'h401615400401407E0402507D42D0507D42C019000B0040160B01541640F04016;
defparam ram_1024_x_18.INIT_08  = 256'h42B0510442A05098429050D14280A2F01210119054165DF04D02AF0F1F90AAFB;
defparam ram_1024_x_18.INIT_09  = 256'h880150A0483CF680C614C7F950D147004016510142E050FF42D0510442C050EB;
defparam ram_1024_x_18.INIT_0A  = 256'h5CB19FE04E041FD0CFFA01051FD050AA2F801FD05CA79FE04E031FD0CDFE1D60;
defparam ram_1024_x_18.INIT_0B  = 256'hCFFC01051FD050BE2F801FD05CBB9FE04E051FD0CFFB01051FD050B42F801FD0;
defparam ram_1024_x_18.INIT_0C  = 256'hCFF80F01CFF80F0050164700CFFD01051FD050C82F801FD05CC59FE04E061FD0;
defparam ram_1024_x_18.INIT_0D  = 256'hFFD07FE08E0150E45D801DE054E25F607FE00E0050E8C80150E84800C6144016;
defparam ram_1024_x_18.INIT_0E  = 256'h46404016C7F354EF46014016CFF80F0040A288017D80C80140D78E0140DB8D01;
defparam ram_1024_x_18.INIT_0F  = 256'hC7F040E808005416467B4016C7F554FB46114016C7F454F746104016C7F754F3;
defparam ram_1024_x_18.INIT_10  = 256'hDFE00E060E060E060E068F0C41068E01590ACF0C0E0040164016C6F2C7F14016;
defparam ram_1024_x_18.INIT_11  = 256'h018005610180054D01800565018005740180056101800547014D0510016AA000;
defparam ram_1024_x_18.INIT_12  = 256'h014D05200180055D018005740180055B01800520018005490180052D0180056E;
defparam ram_1024_x_18.INIT_13  = 256'h0180056501800576018005610180057201800547018005200180052E01800553;
defparam ram_1024_x_18.INIT_14  = 256'hA50F51532510A0000180057401800573018005720180056F018005680180056E;
defparam ram_1024_x_18.INIT_15  = 256'h040604060407145001970166C408A4F01450A0000157C5C0A50FA0000157C580;
defparam ram_1024_x_18.INIT_16  = 256'h01A0016601A50166043001A5A0000191C490A4F8A000C49004F0019B01660406;
defparam ram_1024_x_18.INIT_17  = 256'hA00001A001A0015705010157050C0157050601570528019B01660420019B0166;
defparam ram_1024_x_18.INIT_18  = 256'hC49004F0019B0191C4900406040604070407145001970191C490C40CA4F01450;
defparam ram_1024_x_18.INIT_19  = 256'hA000559CC10101970128A0005598C001000BA000C490E4010197C490E401A000;
defparam ram_1024_x_18.INIT_1A  = 256'h4C00A00055ABC40101A50432A00055A6C30101A00314A00055A1C201019B0219;
defparam ram_1024_x_18.INIT_1B  = 256'h000000008001AA3FCA02EC3F4C0851BC2A80CA01EC3E4C0151B72A40DAC0ACC0;
defparam ram_1024_x_18.INIT_1C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_1F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_20  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_21  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_22  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_23  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_24  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_25  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_26  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_27  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_28  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_29  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_2F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_30  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_31  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_32  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_33  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_34  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_35  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_36  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_37  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_38  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_39  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INIT_3F  = 256'h41AF000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_00 = 256'hC337433737403030D3683DD378C38334CD334F777777777430DDDE22AA00000B;
defparam ram_1024_x_18.INITP_01 = 256'hB37B7B7B7B78D1DD874D0DD788DB34D0B34D0B34D0B34D08766DF77777740D00;
defparam ram_1024_x_18.INITP_02 = 256'hBF3333CFFF3B8A3EA8F02C2C36CCCCCCCCCCCCCCCCCCCCCCCCCCCCCE2A9DD3EB;
defparam ram_1024_x_18.INITP_03 = 256'h000000000000000000000000000000000C2348D02DCB72DCB72D28E28FAA8F80;
defparam ram_1024_x_18.INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_1024_x_18.INITP_07 = 256'hC000000000000000000000000000000000000000000000000000000000000000;
  BSCAN_SPARTAN3 v2_bscan(   
       .TDO1(tdo1),
       .TDO2(tdo2),
            .UPDATE(update),
             .SHIFT(shift),
             .RESET(reset),
               .TDI(tdi),
              .SEL1(sel1),
             .DRCK1(drck1),
              .SEL2(sel2),
             .DRCK2(drck2),
    .CAPTURE(capture));
    
  //buffer signal used as a clock
  BUFG upload_clock(
          .I(drck1),
          .O(drck1_buf));
  // Assign the reset to be active whenever the uploading subsystem is active
  assign proc_reset = sel1;
  defparam srlC1.INIT = 16'h0000;
  SRLC16E srlC1 (   
              .D(tdi),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[10]),
            .Q15(jaddr[8]));
            
  FD flop1(
             .D(jaddr[10]),
             .Q(jaddr[9]),
             .C(drck1_buf));
  defparam srlC2.INIT = 16'h0000;
  SRLC16E srlC2 (   
              .D(jaddr[8]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[7]),
            .Q15(tap5));
            
  FD flop2 ( 
             .D(jaddr[7]),
             .Q(jaddr[6]),
             .C(drck1_buf));
  defparam srlC3.INIT = 16'h0000;
  SRLC16E srlC3(   
              .D(tap5),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[5]),
            .Q15(jaddr[3]));
  
  FD flop3 ( 
             .D(jaddr[5]),
             .Q(jaddr[4]),
             .C(drck1_buf));
  defparam srlC4.INIT = 16'h0000;
  SRLC16E srlC4 (   
              .D(jaddr[3]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[2]),
            .Q15(tap11));
  
  FD flop4 ( 
             .D(jaddr[2]),
             .Q(jaddr[1]),
             .C(drck1_buf));
  defparam srlC5.INIT = 16'h0000;
  SRLC16E srlC5 (   
              .D(tap11),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jaddr[0]),
            .Q15(jdata[7]));
            
  FD flop5 ( 
             .D(jaddr[0]),
             .Q(jparity[0]),
             .C(drck1_buf));
  defparam srlC6.INIT = 16'h0000;
    SRLC16E srlC6(   
             .D(jdata[7]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[6]),
            .Q15(tap17));
  
  FD flop6 ( 
             .D(jdata[6]),
             .Q(jdata[5]),
             .C(drck1_buf));
  defparam srlC7.INIT = 16'h0000;
  SRLC16E srlC7 (   
              .D(tap17),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[4]),
            .Q15(jdata[2]));
  
  FD flop7 ( 
             .D(jdata[4]),
             .Q(jdata[3]),
             .C(drck1_buf));
  defparam srlC8.INIT = 16'h0000;
  SRLC16E srlC8 (   
             .D(jdata[2]),
             .CE(1'b1),
            .CLK(drck1_buf),
             .A0(1'b1),
             .A1(1'b0),
             .A2(1'b1),
             .A3(1'b1),
              .Q(jdata[1]),
            .Q15(tdo1));
  FD flop8 ( 
             .D(jdata[1]),
             .Q(jdata[0]),
             .C(drck1_buf));
endmodule
